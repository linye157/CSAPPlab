module count6_tb(

    );
    reg rst;
    reg clk;
    reg en;
    wire [2:0] count;
    wire co;
    initial begin
        rst = 0;
        clk = 0;
        en = 0;
        #100
        rst = 1;
        #40
        rst = 0;
        en = 1;
    end
    
    always #10 clk = ~clk;
    count_6 count6(rst,clk,en,count,co);    
endmodule